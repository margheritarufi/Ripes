//These are parameters that the designer can change

`define TGDI_WIDTH 1
`define TGDO_WIDTH 1
`define TGA_WIDTH 1
`define TGC_WIDTH 1
`define SEL_WIDTH 1
